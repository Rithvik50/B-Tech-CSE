module not2(b, a);
input a;
output b;
assign b = !a;
endmodule